MACRO LATCH
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN LATCH 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal1 ;
        RECT 0.00000000 30500.00000000 56000.00000000 33500.00000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal1 ;
        RECT 0.00000000 -1500.00000000 56000.00000000 1500.00000000 ;
    END
  END GND

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 27000.00000000 9500.00000000 29000.00000000 19500.00000000 ;
    END
  END CLK

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 15000.00000000 13500.00000000 17000.00000000 15500.00000000 ;
    END
  END D

  PIN Q
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 39000.00000000 13500.00000000 41000.00000000 15500.00000000 ;
    END
  END Q


END LATCH
